//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Roseek Ltd. All rights reserved
// -----------------------------------------------------------------------------
// FILE NAME : 
// DEPARTMENT : FPGA team
// AUTHOR : Sha Craig
// AUTHOR'S EMAIL : 
// -----------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION  DATE            AUTHOR      DESCRIPTION
// 0.1      2016-05-30      Craig       Creat
//----------------------------------------------------------------------------- 
// REUSE ISSUES
// Reset Strategy : None
// Clock Domains :
// Critical Timing :
// Test Features :
// Asynchronous I/F :
// Scan Methodology :
// Instantiations :
// Synthesizable : Y
// Other :
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ps / 1ps

module mt9v034_bridge #(
parameter TCQ = 100,
parameter SIM = 1)(
input rst,

input dlck_p,
input dlck_n,
input dlo_p,
input dlo_n,

input im_oe,
output mmcm_locked,
output align_err,

output pixel_clk,
output im_vsync,
output im_hsync,
output im_valid,
output[15: 0] im_dout
);

genvar i;

/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/


/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/
wire dlo_clk;
wire dlo_valid;
wire[17: 0] dlo;

wire dlo_align_valid;
wire[17: 0] dlo_align;

(* MARK_DEBUG = "TRUE" *)
wire im_vsync_i;
(* MARK_DEBUG = "TRUE" *)
wire im_hsync_i;
(* MARK_DEBUG = "TRUE" *)
wire im_valid_i;
(* MARK_DEBUG = "TRUE" *)
wire[15: 0] im_data_i;


/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
(* ASYNC_REG = "TRUE" *)
reg[3 : 0] im_oe_sync = 4'H0;
reg im_oe_d = 1'B0;

reg im_vsync_d;
reg im_hsync_d;
reg im_valid_d;
reg[15: 0] im_dout_d;

reg im_vsync_dd;
reg im_hsync_dd;
reg im_valid_dd;
reg[15: 0] im_dout_dd;

/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/**************************************  Start instants Declaration  ***************************************/
/***********************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : instance
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
mt9v034_lvds_iserdes #(
.TCQ( TCQ),
.SIM( SIM))
mt9v034_lvds_iserdes_inst(
.rst( rst),

.dlck_p( dlck_p),
.dlck_n( dlck_n),
.dlo_p( dlo_p),
.dlo_n( dlo_n),

.mmcm_locked( mmcm_locked),
.pixel_clk( pixel_clk),
.dlo_clk( dlo_clk),
.dlo_valid( dlo_valid),
.dlo( dlo)
);


//------------------------------------------------------------------------------
// NAME : 
// TYPE : instance
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
mt9v034_lvds_bit_align #(
.TCQ( TCQ),
.SIM( SIM))
mt9v034_lvds_bit_align_inst(
.rst( rst),

.dlo_clk( dlo_clk),
.dlo_valid_i( dlo_valid),
.dlo_i( dlo),

.align_err( align_err),
.dlo_valid_o( dlo_align_valid),
.dlo_o( dlo_align)
);

//------------------------------------------------------------------------------
// NAME : 
// TYPE : instance
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
mt9v034_lvds_protocol_decode #(
.TCQ( TCQ),
.SIM( SIM))
mt9v034_lvds_protocol_decode_inst(
.rst( rst),

.dlo_clk( dlo_clk),
.dlo_valid_i( dlo_align_valid),
.dlo_i( dlo_align),

.im_vsync( im_vsync_i),
.im_hsync( im_hsync_i),
.im_valid( im_valid_i),
.im_data( im_data_i)
);



/*************************************************************************************************************/
/***************************************  End of instants Declaration  ***************************************/
/*************************************************************************************************************/


/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge pixel_clk or negedge im_oe)
begin
    if( ~im_oe) begin
        im_oe_sync <= #TCQ 4'H0;
    end else begin
        im_oe_sync <= #TCQ { im_oe_sync[2 : 0], 1'B1};
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge pixel_clk)
begin
    if( ~im_oe_sync[ 3]) begin
        im_oe_d <= #TCQ 1'B0;
    end else begin
        if( im_vsync_i) begin
            im_oe_d <= #TCQ 1'B1;
        end else begin
            im_oe_d <= #TCQ im_oe_d;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge pixel_clk)
begin
    im_vsync_d <= #TCQ im_vsync_i;
    im_hsync_d <= #TCQ im_hsync_i;
    im_valid_d <= #TCQ im_valid_i;

    if( im_oe_d) begin
        im_vsync_dd <= #TCQ im_vsync_d;
        im_hsync_dd <= #TCQ im_hsync_d;
        im_valid_dd <= #TCQ im_valid_d;
    end else begin
        im_vsync_dd <= #TCQ 1'B1;
        im_hsync_dd <= #TCQ 1'B1;
        im_valid_dd <= #TCQ 1'B0;
    end

    im_dout_d <= #TCQ im_dout_i;
    im_dout_dd <= #TCQ im_dout_d;
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : assignment
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
assign im_vsync = im_vsync_dd;
assign im_hsync = im_hsync_dd;
assign im_valid = im_valid_dd;
assign im_dout = im_dout_dd;

/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/






/*************************************************************************************************************/
/*********************************  Begin simulation information display  ************************************/
/*************************************************************************************************************/
// synthesis translate_off


// synthesis translate_on
/*************************************************************************************************************/
/*********************************  End simulation information display  **************************************/
/*************************************************************************************************************/
endmodule
