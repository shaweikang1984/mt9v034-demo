//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Roseek Ltd. All rights reserved
// -----------------------------------------------------------------------------
// FILE NAME : 
// DEPARTMENT : FPGA team
// AUTHOR : Sha Craig
// AUTHOR'S EMAIL : 
// -----------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION  DATE            AUTHOR      DESCRIPTION
// 0.1      2016-05-30      Craig       Creat
//----------------------------------------------------------------------------- 
// REUSE ISSUES
// Reset Strategy : None
// Clock Domains :
// Critical Timing :
// Test Features :
// Asynchronous I/F :
// Scan Methodology :
// Instantiations :
// Synthesizable : Y
// Other :
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ps / 1ps

module mt9v034_lvds_bit_align #(
parameter TCQ = 100,
parameter SIM = 1)(
input rst,

input dlo_clk,

input dlo_valid_i,
input[17: 0] dlo_i,

output align_err,
output dlo_valid_o,
output[17: 0] dlo_o
);

genvar i;
genvar j;
/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/

localparam C_IDLE = 0;
localparam C_DECT = 1;
localparam C_BSLIP = 2;
localparam C_HOLD = 3;
localparam C_ALIGNED = 4;
localparam C_ERROR = 5;
/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/
wire rst_i;

wire frame_valid;

wire[35: 0] dlo_align_package_l;
wire[35: 0] dlo_align_package_h;


/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
(* ASYNC_REG = "TRUE" *)
reg[7 : 0] rst_sync = 8'Hff;

reg dlo_valid_d = 1'B0;
reg dlo_valid_dd = 1'B0;

reg[17: 0] dlo_d = 18'D0;
reg[17: 0] dlo_dd = 18'D0;

reg[17: 0] align_shift = 18'D1;

reg[5 : 0] align_cs = 6'B00_0001;
reg[5 : 0] align_ns;

reg[11: 0] frame_valid_cnt = 12'D0;

reg[17: 0] dlo_align = 18'D0;
/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/**************************************  Start instants Declaration  ***************************************/
/***********************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : instance
// -----------------------------------------------------------------------------
// PURPOSE : srl implement by dsp
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
dlo_srl dlo_srl_inst_h(
.CLK( dlo_clk), // input wire CLK
.A( align_shift), // input wire [17 : 0] A
.B( dlo_dd), // input wire [17 : 0] B
.P( dlo_align_package_h) // output wire [35 : 0] P
);

//------------------------------------------------------------------------------
// NAME : 
// TYPE : instance
// -----------------------------------------------------------------------------
// PURPOSE : srl implement by dsp
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
dlo_srl dlo_srl_inst_l(
.CLK( dlo_clk), // input wire CLK
.A( align_shift), // input wire [17 : 0] A
.B( dlo_d), // input wire [17 : 0] B
.P( dlo_align_package_l) // output wire [35 : 0] P
);

/*************************************************************************************************************/
/***************************************  End of instants Declaration  ***************************************/
/*************************************************************************************************************/


/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/

/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk or posedge rst)
begin
      if( rst) begin
            rst_sync <= #TCQ 8'Hff;
      end else begin
            rst_sync <= #TCQ { rst_sync[6 : 0], 1'B0};
      end
end

assign rst_i = rst_sync[ 31];

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk)
begin
    dlo_d <= #TCQ dlo_i;
    dlo_dd <= #TCQ dlo_d;

    dlo_valid_d <= #TCQ dlo_valid_i;
    dlo_valid_dd <= #TCQ dlo_valid_d;
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk)
begin
    dlo_align <= #TCQ dlo_align_package_h[17: 0] | dlo_align_package_l[35:18];
end

assign frame_valid = ( ~dlo_align[ 17]) & ( dlo_align[ 0]);

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk or posedge rst_i)
begin
    if( rst_i) begin
        align_cs[ C_IDLE] <= #TCQ 1'B1;
        align_cs[ C_DECT] <= #TCQ 1'B0;
        align_cs[ C_BSLIP] <= #TCQ 1'B0;
        align_cs[ C_HOLD] <= #TCQ 1'B0;
        align_cs[ C_ALIGNED] <= #TCQ 1'B0;
        align_cs[ C_ERROR] <= #TCQ 1'B0;
    end else begin
        align_cs <= #TCQ align_ns;
    end
end

always @*
begin
    align_ns = 'D0;

    case( 1'B1)
        align_cs[ C_IDLE]:      begin
                                    if( dlo_valid_dd) begin
                                        align_ns[ C_DECT] = 1'B1;
                                    end
                                end
        align_cs[ C_DECT]:      begin
                                    if( ~frame_valid) begin
                                        align_ns[ C_BSLIP] = 1'B1;
                                    end else begin
                                        if( &frame_valid_cnt) begin
                                            align_ns[ C_ALIGNED] = 1'B1;
                                        end else begin
                                            align_ns[ C_DECT] = 1'B1;
                                        end
                                    end
                                end
        align_cs[ C_BSLIP]:     begin
                                    if( align_shift[ 0]) begin
                                        align_ns[ C_ERROR] = 1'B1;
                                    end else begin
                                        align_ns[ C_HOLD] = 1'B1;
                                    end
                                end
        align_cs[ C_HOLD]:      begin
                                    align_ns[ C_DECT] = 1'B1;
                                end
        align_cs[ C_ALIGNED]:   begin
                                    if( ~frame_valid) begin
                                        align_ns[ C_ERROR] = 1'B1;
                                    end else begin
                                        align_ns[ C_ALIGNED] = 1'B1;
                                    end
                                end
        align_cs[ C_ERROR]:     begin
                                    align_ns[ C_ERROR] = 1'B1;
                                end
    endcase
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk)
begin
    if( align_ns[ C_IDLE]) begin
        align_shift <= #TCQ 18'D1;
    end else if( align_ns[ C_BSLIP]) begin
        align_shift <= #TCQ { align_shift[16: 0], align_shift[ 17]};
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk)
begin
    if( align_cs[ C_DECT] & frame_valid) begin
        frame_valid_cnt <= #TCQ frame_valid_cnt + 1'B1;
    end else begin
        frame_valid_cnt <= 12'D0;
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : assignment
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
assign dlo_o = dlo_align;
assign dlo_valid_o = align_cs[ C_ALIGNED];

assign align_err = align_cs[ C_ERROR];

/*************************************************************************************************************/
/*********************************  Begin simulation information display  ************************************/
/*************************************************************************************************************/
// synthesis translate_off


// synthesis translate_on
/*************************************************************************************************************/
/*********************************  End simulation information display  **************************************/
/*************************************************************************************************************/
endmodule
