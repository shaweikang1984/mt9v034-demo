//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Roseek Ltd. All rights reserved
// -----------------------------------------------------------------------------
// FILE NAME : 
// DEPARTMENT : FPGA team
// AUTHOR : Sha Craig
// AUTHOR'S EMAIL : 
// -----------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION  DATE            AUTHOR      DESCRIPTION
// 0.1      2016-05-30      Craig       Creat
//----------------------------------------------------------------------------- 
// REUSE ISSUES
// Reset Strategy : None
// Clock Domains :
// Critical Timing :
// Test Features :
// Asynchronous I/F :
// Scan Methodology :
// Instantiations :
// Synthesizable : Y
// Other :
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ps / 1ps

module mt9v034_lvds_protocol_decode #(
parameter TCQ = 100,
parameter SIM = 1)(
input rst,

input dlo_clk,
input dlo_valid_i,
input[17: 0] dlo_i,

output im_vsync,
output im_hsync,
output im_valid,
output[15: 0] im_data
);

genvar i;
genvar j;
/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/

localparam fsav = 8'H0;
localparam feav = 8'H3;
localparam sav = 8'H1;
localparam eav = 8'H2;

/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/
wire rst_i;

/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/

/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
(* ASYNC_REG = "TRUE" *)
reg[3: 0] rst_sync = 4'Hf;

reg im_vsync_d = 1'B1;
reg im_hsync_d = 1'B1;

/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/**************************************  Start instants Declaration  ***************************************/
/***********************************************************************************************************/


/*************************************************************************************************************/
/***************************************  End of instants Declaration  ***************************************/
/*************************************************************************************************************/


/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk or posedge rst)
begin
      if( rst) begin
            rst_sync <= #TCQ 4'Hf;
      end else begin
            rst_sync <= #TCQ { rst_sync[2 : 0], 1'B0};
      end
end

assign rst_i = rst_sync[ 3];

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk or posedge rst)
begin
    if( rst) begin
        im_vsync_d <= #TCQ 1'B1;
    end else if( dlo_valid_i) begin
        if( dlo_i[8 : 1] == fsav) begin
            im_vsync_d <= #TCQ 1'B0;
        end else if( dlo_i[8 : 1] == feav) begin
            im_vsync_d <= #TCQ 1'B0;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge dlo_clk or posedge rst)
begin
    if( rst) begin
        im_hsync_d <= #TCQ 1'B1;
    end else if( dlo_valid_i) begin
        if( dlo_i[8 : 1] == sav) begin
            im_hsync_d <= #TCQ 1'B0;
        end else if( dlo_i[8 : 1] == eav) begin
            im_hsync_d <= #TCQ 1'B0;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : assignment
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
assign im_vsync = im_vsync_d;
assign im_hsync = im_hsync_d;
assign im_valid = ~im_hsync_d;
assign im_data = dlo_i[16: 1];


/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/






/*************************************************************************************************************/
/*********************************  Begin simulation information display  ************************************/
/*************************************************************************************************************/
// synthesis translate_off


// synthesis translate_on
/*************************************************************************************************************/
/*********************************  End simulation information display  **************************************/
/*************************************************************************************************************/
endmodule
