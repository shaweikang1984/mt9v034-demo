`define test