//////////////////////////////////////////////////////////////////////////////////
// Copyright (c) Roseek Ltd. All rights reserved
// -----------------------------------------------------------------------------
// FILE NAME : 
// DEPARTMENT : FPGA team
// AUTHOR : Sha Craig
// AUTHOR鈥橲 EMAIL : shaweikang@roseek.com
// -----------------------------------------------------------------------------
// RELEASE HISTORY
// VERSION  DATE            AUTHOR      DESCRIPTION
// 0.1      2014-12-03      Craig       Creat
//----------------------------------------------------------------------------- 
// REUSE ISSUES
// Reset Strategy : None
// Clock Domains :
// Critical Timing :
// Test Features :
// Asynchronous I/F :
// Scan Methodology :
// Instantiations :
// Synthesizable : Y
// Other :
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ps / 1ps

module mt9v034_i2c_if #(
parameter TCQ = 100,
parameter SIM = 0)(
input rst,
input clk,

input trans_trg,
input[3 : 0] trans_bit_num,
input[10: 0] trans_din,
output[9 : 0] trans_dout,
output trans_done,

output scl_oen,
output scl_o,
input scl_i,
output sda_oen,
output sda_o,
input sda_i
);


/***********************************************************************************************************/
/*************************************  Start Parameter Declaration  ***************************************/
/***********************************************************************************************************/
localparam T_IDLE = 0;
localparam T_START = 1;
localparam T_TRANS = 2;
localparam T_STOP = 3;
localparam T_DONE = 4;
/***********************************************************************************************************/
/***************************************  End Parameter Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/******************************************  Start Wire Declaration  ***************************************/
/***********************************************************************************************************/
wire rst_i;
/*************************************************************************************************************/
/*****************************************  End Wire Declaration  ********************************************/
/*************************************************************************************************************/



/***********************************************************************************************************/
/*************************************  Start Registers Declaration  ***************************************/
/***********************************************************************************************************/
(* ASYNC_REG = "true" *)
reg[3 : 0] rst_sync = 4'Hf;

(* ASYNC_REG = "true" *)
reg scl_i_d0 = 1'B1;
(* ASYNC_REG = "true" *)
reg scl_i_d1 = 1'B1;
reg scl_i_d2 = 1'B1;
reg scl_i_d3 = 1'B1;
reg scl_i_neg = 1'B0;
reg scl_i_pos = 1'B0;

(* ASYNC_REG = "true" *)
reg sda_i_d0 = 1'B1;
(* ASYNC_REG = "true" *)
reg sda_i_d1 = 1'B1;

reg[9 : 0] clk_div_cnt = 10'D0;
reg clk_div_en = 1'B0;

(* fsm_encoding = "one-hot" *)
reg[4 : 0] t_cs = 5'B0_0001;
reg[4 : 0] t_ns;

reg trans_done_d = 1'B0;

reg[3 : 0] trans_cnt = 4'D0;
reg[10: 0] trans_srl = 11'B111_1111_1111;

reg[9 : 0] reseive_srl = 10'D0;

reg sda_oen_d = 1'B1;
reg sda_oen_dd = 1'B1;
reg sda_oen_ddd = 1'B1;
reg sda_oen_dddd = 1'B1;
reg sda_oen_ddddd = 1'B1;
reg sda_oen_dddddd = 1'B1;
reg scl_oen_d = 1'B1;

/***********************************************************************************************************/
/***************************************  End Registers Declaration  ***************************************/
/***********************************************************************************************************/

/***********************************************************************************************************/
/*****************************************  Start instances Declaration  ************************************/
/***********************************************************************************************************/
//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst)
begin
    if( rst) begin
        rst_sync <= #TCQ 4'H0;
    end else begin
        rst_sync <= #TCQ { rst_sync[2 : 0], 1'B0};
    end
end

assign rst_i = rst_sync[ 3];


//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk)
begin
    scl_i_d0 <= #TCQ scl_i;
    scl_i_d1 <= #TCQ scl_i_d0;
    scl_i_d2 <= #TCQ scl_i_d1;
    scl_i_d3 <= #TCQ scl_i_d2;
    scl_i_neg <= #TCQ scl_i_d3 & ( ~scl_i_d2);
    scl_i_pos <= #TCQ scl_i_d2 & ( ~scl_i_d3);
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk)
begin
    sda_i_d0 <= #TCQ sda_i;
    sda_i_d1 <= #TCQ sda_i_d0;
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : fsm
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        t_cs[ T_IDLE] <= #TCQ 1'B1;
        t_cs[ T_START] <= #TCQ 1'B0;
        t_cs[ T_TRANS] <= #TCQ 1'B0;
        t_cs[ T_STOP] <= #TCQ 1'B0;
        t_cs[ T_DONE] <= #TCQ 1'B0;
    end else begin
        t_cs <= #TCQ t_ns;
    end
end

always @*
begin
    t_ns = 'D0;

    (* full_case, parallel_case *)
    case( 1'B1)
        t_cs[ T_IDLE]:  begin
                            if( trans_trg) begin
                                t_ns[ T_START] = 1'B1;
                            end else begin
                                t_ns[ T_IDLE] = 1'B1;
                            end
                        end
        t_cs[ T_START]: begin
                            if( clk_div_en) begin
                                t_ns[ T_TRANS] = 1'B1;
                            end else begin
                                t_ns[ T_START] = 1'B1;
                            end
                        end
        t_cs[ T_TRANS]: begin
                            if( trans_cnt == 4'D0) begin
                                t_ns[ T_STOP] = 1'B1;
                            end else begin
                                t_ns[ T_TRANS] = 1'B1;
                            end
                        end
        t_cs[ T_STOP]:  begin
                            if( clk_div_en) begin
                                t_ns[ T_DONE] = 1'B1;
                            end else begin
                                t_ns[ T_STOP] = 1'B1;
                            end
                        end
        t_cs[ T_DONE]:  begin
                            if( clk_div_en) begin
                                t_ns[ T_IDLE] = 1'B1;
                            end else begin
                                t_ns[ T_DONE] = 1'B1;
                            end
                        end
    endcase
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        { clk_div_en, clk_div_cnt} <= #TCQ 'D0;
    end else begin
        if( t_ns[ T_IDLE]) begin
            { clk_div_en, clk_div_cnt} <= #TCQ 'D0;
        end else begin
            { clk_div_en, clk_div_cnt} <= #TCQ clk_div_cnt + 1'B1;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        trans_cnt <= #TCQ 4'D0;
    end else begin
        if( trans_trg) begin
            trans_cnt <= #TCQ trans_bit_num;
        end else if( clk_div_en & ( ~scl_oen_d)) begin
            trans_cnt <= #TCQ trans_cnt - 1'B1;
        end else begin
            trans_cnt <= #TCQ trans_cnt;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk)
begin
    if( trans_trg) begin
        trans_srl <= #TCQ { trans_din[ 10], // start bit
                            trans_din[9 : 2],
                            trans_din[ 1], // ack bit
                            trans_din[ 0]}; // stop bit
    end else if( scl_i_neg) begin
        trans_srl <= #TCQ { trans_srl[9 : 0], 1'B0};
    end else begin
        trans_srl <= #TCQ trans_srl;
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk)
begin
    if( trans_trg) begin
        reseive_srl <= #TCQ 10'D0;
    end else if( scl_i_pos) begin
        reseive_srl <= #TCQ { reseive_srl[8 : 0], sda_i_d1};
    end
end


assign trans_dout = reseive_srl;
//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        sda_oen_d <= #TCQ 1'B1;
    end else begin
        (* full_case, parallel_case *)
        case( 1'B1)
            t_ns[ T_IDLE]:  begin
                                sda_oen_d <= #TCQ 1'B1;
                            end
            t_ns[ T_START]: begin // i2c start bit
                                sda_oen_d <= #TCQ trans_srl[ 10];
                            end
            t_ns[ T_TRANS]: begin // i2c data
                                sda_oen_d <= #TCQ trans_srl[ 10];
                            end
            t_ns[ T_STOP]:  begin // i2c stop bit
                                sda_oen_d <= #TCQ trans_srl[ 10];
                            end
            t_ns[ T_DONE]:  begin
                                sda_oen_d <= #TCQ 1'B1;
                            end
        endcase
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        scl_oen_d <= #TCQ 1'B1;
    end else begin
        (* full_case, parallel_case *)
        case( 1'B1)
            t_ns[ T_IDLE]:  begin
                                scl_oen_d <= #TCQ 1'B1;
                            end
            t_ns[ T_DONE]:  begin
                                scl_oen_d <= #TCQ 1'B1; 
                            end
            default:        begin
                                if( clk_div_en) begin
                                    scl_oen_d <= #TCQ ~scl_oen_d;
                                end else begin
                                    scl_oen_d <= #TCQ scl_oen_d;
                                end
                            end
        endcase
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk or posedge rst_i)
begin
    if( rst_i) begin
        trans_done_d <= #TCQ 1'B1;
    end else begin
        if( trans_trg) begin
            trans_done_d <= #TCQ 1'B0;
        end else if( t_cs[ T_DONE] & clk_div_en) begin
            trans_done_d <= #TCQ 1'B1;
        end else begin
            trans_done_d <= #TCQ trans_done_d;
        end
    end
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : assignment
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
assign trans_done = trans_done_d;


//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
always @( posedge clk)
begin
    sda_oen_dd <= #TCQ sda_oen_d;
    sda_oen_ddd <= #TCQ sda_oen_dd;
    sda_oen_dddd <= #TCQ sda_oen_ddd;
    sda_oen_ddddd <= #TCQ sda_oen_dddd;
    sda_oen_dddddd <= #TCQ sda_oen_ddddd;
end

//------------------------------------------------------------------------------
// NAME : 
// TYPE : assignment
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------
assign scl_oen = scl_oen_d;
assign scl_o = 1'B0;

assign sda_oen = sda_oen_dddddd;
assign sda_o = 1'B0;
/***********************************************************************************************************/
/****************************************  End of instants Declaration  ************************************/
/***********************************************************************************************************/


/*************************************************************************************************************/
/*********************************  Start Design RTL Description  ********************************************/
/*************************************************************************************************************/

//------------------------------------------------------------------------------
// NAME : 
// TYPE : process
// -----------------------------------------------------------------------------
// PURPOSE : 
// -----------------------------------------------------------------------------
// Other : 
//------------------------------------------------------------------------------

/*************************************************************************************************************/
/***********************************  End Design RTL Description  ********************************************/
/*************************************************************************************************************/



/*************************************************************************************************************/
/*********************************  Begin simulation information display  ************************************/
/*************************************************************************************************************/
// synthesis translate_off


// synthesis translate_on
/*************************************************************************************************************/
/*********************************  End simulation information display  **************************************/
/*************************************************************************************************************/
endmodule
